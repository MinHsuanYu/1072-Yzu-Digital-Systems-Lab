module lab6(SW,LED);
	input [9:0]SW;
	output [9:0]LED;
	assign LED = SW;
endmodule 