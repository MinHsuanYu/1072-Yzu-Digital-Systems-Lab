library verilog;
use verilog.vl_types.all;
entity S1061534_lab5_test is
end S1061534_lab5_test;
